   // NESCTRL
   input             nesctrl_ctrl1_q7,
   input             nesctrl_ctrl2_q7,
   output            nesctrl_pl1,
   output            nesctrl_pl2,
   output            nesctrl_clk1,
   output            nesctrl_clk2,
   output [8-1:0]    nesctrl_ctrl2_data,
