   // NESCTRL
   input             nesctrl_ctrl1_q7,
   input             nesctrl_ctrl2_q7,
   output            nesctrl_pl,
   output [16-1:0]   nesctrl_ctrl1_data,
   output [16-1:0]   nesctrl_ctrl2_data,
